`include "fa.v"
`include "ha.v"
`include "cp_acc.v"
`include "cp_app.v"
module wallace_acc(a,b,sum);
	input[15:0] a,b;
  

	output[31:0] sum;
  
	wire ground_z;
	assign ground_z = 1'b0;
	//-------------------------------------------AND layer---------------------------------------//
	wire P_0_0;
	wire P_0_1;
	wire P_0_2;
	wire P_0_3;
	wire P_0_4;
	wire P_0_5;
	wire P_0_6;
	wire P_0_7;
	wire P_0_8;
	wire P_0_9;
	wire P_0_10;
	wire P_0_11;
	wire P_0_12;
	wire P_0_13;
	wire P_0_14;
	wire P_0_15;
	wire P_1_0;
	wire P_1_1;
	wire P_1_2;
	wire P_1_3;
	wire P_1_4;
	wire P_1_5;
	wire P_1_6;
	wire P_1_7;
	wire P_1_8;
	wire P_1_9;
	wire P_1_10;
	wire P_1_11;
	wire P_1_12;
	wire P_1_13;
	wire P_1_14;
	wire P_1_15;
	wire P_2_0;
	wire P_2_1;
	wire P_2_2;
	wire P_2_3;
	wire P_2_4;
	wire P_2_5;
	wire P_2_6;
	wire P_2_7;
	wire P_2_8;
	wire P_2_9;
	wire P_2_10;
	wire P_2_11;
	wire P_2_12;
	wire P_2_13;
	wire P_2_14;
	wire P_2_15;
	wire P_3_0;
	wire P_3_1;
	wire P_3_2;
	wire P_3_3;
	wire P_3_4;
	wire P_3_5;
	wire P_3_6;
	wire P_3_7;
	wire P_3_8;
	wire P_3_9;
	wire P_3_10;
	wire P_3_11;
	wire P_3_12;
	wire P_3_13;
	wire P_3_14;
	wire P_3_15;
	wire P_4_0;
	wire P_4_1;
	wire P_4_2;
	wire P_4_3;
	wire P_4_4;
	wire P_4_5;
	wire P_4_6;
	wire P_4_7;
	wire P_4_8;
	wire P_4_9;
	wire P_4_10;
	wire P_4_11;
	wire P_4_12;
	wire P_4_13;
	wire P_4_14;
	wire P_4_15;
	wire P_5_0;
	wire P_5_1;
	wire P_5_2;
	wire P_5_3;
	wire P_5_4;
	wire P_5_5;
	wire P_5_6;
	wire P_5_7;
	wire P_5_8;
	wire P_5_9;
	wire P_5_10;
	wire P_5_11;
	wire P_5_12;
	wire P_5_13;
	wire P_5_14;
	wire P_5_15;
	wire P_6_0;
	wire P_6_1;
	wire P_6_2;
	wire P_6_3;
	wire P_6_4;
	wire P_6_5;
	wire P_6_6;
	wire P_6_7;
	wire P_6_8;
	wire P_6_9;
	wire P_6_10;
	wire P_6_11;
	wire P_6_12;
	wire P_6_13;
	wire P_6_14;
	wire P_6_15;
	wire P_7_0;
	wire P_7_1;
	wire P_7_2;
	wire P_7_3;
	wire P_7_4;
	wire P_7_5;
	wire P_7_6;
	wire P_7_7;
	wire P_7_8;
	wire P_7_9;
	wire P_7_10;
	wire P_7_11;
	wire P_7_12;
	wire P_7_13;
	wire P_7_14;
	wire P_7_15;
	wire P_8_0;
	wire P_8_1;
	wire P_8_2;
	wire P_8_3;
	wire P_8_4;
	wire P_8_5;
	wire P_8_6;
	wire P_8_7;
	wire P_8_8;
	wire P_8_9;
	wire P_8_10;
	wire P_8_11;
	wire P_8_12;
	wire P_8_13;
	wire P_8_14;
	wire P_8_15;
	wire P_9_0;
	wire P_9_1;
	wire P_9_2;
	wire P_9_3;
	wire P_9_4;
	wire P_9_5;
	wire P_9_6;
	wire P_9_7;
	wire P_9_8;
	wire P_9_9;
	wire P_9_10;
	wire P_9_11;
	wire P_9_12;
	wire P_9_13;
	wire P_9_14;
	wire P_9_15;
	wire P_10_0;
	wire P_10_1;
	wire P_10_2;
	wire P_10_3;
	wire P_10_4;
	wire P_10_5;
	wire P_10_6;
	wire P_10_7;
	wire P_10_8;
	wire P_10_9;
	wire P_10_10;
	wire P_10_11;
	wire P_10_12;
	wire P_10_13;
	wire P_10_14;
	wire P_10_15;
	wire P_11_0;
	wire P_11_1;
	wire P_11_2;
	wire P_11_3;
	wire P_11_4;
	wire P_11_5;
	wire P_11_6;
	wire P_11_7;
	wire P_11_8;
	wire P_11_9;
	wire P_11_10;
	wire P_11_11;
	wire P_11_12;
	wire P_11_13;
	wire P_11_14;
	wire P_11_15;
	wire P_12_0;
	wire P_12_1;
	wire P_12_2;
	wire P_12_3;
	wire P_12_4;
	wire P_12_5;
	wire P_12_6;
	wire P_12_7;
	wire P_12_8;
	wire P_12_9;
	wire P_12_10;
	wire P_12_11;
	wire P_12_12;
	wire P_12_13;
	wire P_12_14;
	wire P_12_15;
	wire P_13_0;
	wire P_13_1;
	wire P_13_2;
	wire P_13_3;
	wire P_13_4;
	wire P_13_5;
	wire P_13_6;
	wire P_13_7;
	wire P_13_8;
	wire P_13_9;
	wire P_13_10;
	wire P_13_11;
	wire P_13_12;
	wire P_13_13;
	wire P_13_14;
	wire P_13_15;
	wire P_14_0;
	wire P_14_1;
	wire P_14_2;
	wire P_14_3;
	wire P_14_4;
	wire P_14_5;
	wire P_14_6;
	wire P_14_7;
	wire P_14_8;
	wire P_14_9;
	wire P_14_10;
	wire P_14_11;
	wire P_14_12;
	wire P_14_13;
	wire P_14_14;
	wire P_14_15;
	wire P_15_0;
	wire P_15_1;
	wire P_15_2;
	wire P_15_3;
	wire P_15_4;
	wire P_15_5;
	wire P_15_6;
	wire P_15_7;
	wire P_15_8;
	wire P_15_9;
	wire P_15_10;
	wire P_15_11;
	wire P_15_12;
	wire P_15_13;
	wire P_15_14;
	wire P_15_15;
  
	and A_0_0(P_0_0, a[0], b[0]);
	and A_0_1(P_0_1, a[0], b[1]);
	and A_0_2(P_0_2, a[0], b[2]);
	and A_0_3(P_0_3, a[0], b[3]);
	and A_0_4(P_0_4, a[0], b[4]);
	and A_0_5(P_0_5, a[0], b[5]);
	and A_0_6(P_0_6, a[0], b[6]);
	and A_0_7(P_0_7, a[0], b[7]);
	and A_0_8(P_0_8, a[0], b[8]);
	and A_0_9(P_0_9, a[0], b[9]);
	and A_0_10(P_0_10, a[0], b[10]);
	and A_0_11(P_0_11, a[0], b[11]);
	and A_0_12(P_0_12, a[0], b[12]);
	and A_0_13(P_0_13, a[0], b[13]);
	and A_0_14(P_0_14, a[0], b[14]);
	and A_0_15(P_0_15, a[0], b[15]);
	and A_1_0(P_1_0, a[1], b[0]);
	and A_1_1(P_1_1, a[1], b[1]);
	and A_1_2(P_1_2, a[1], b[2]);
	and A_1_3(P_1_3, a[1], b[3]);
	and A_1_4(P_1_4, a[1], b[4]);
	and A_1_5(P_1_5, a[1], b[5]);
	and A_1_6(P_1_6, a[1], b[6]);
	and A_1_7(P_1_7, a[1], b[7]);
	and A_1_8(P_1_8, a[1], b[8]);
	and A_1_9(P_1_9, a[1], b[9]);
	and A_1_10(P_1_10, a[1], b[10]);
	and A_1_11(P_1_11, a[1], b[11]);
	and A_1_12(P_1_12, a[1], b[12]);
	and A_1_13(P_1_13, a[1], b[13]);
	and A_1_14(P_1_14, a[1], b[14]);
	and A_1_15(P_1_15, a[1], b[15]);
	and A_2_0(P_2_0, a[2], b[0]);
	and A_2_1(P_2_1, a[2], b[1]);
	and A_2_2(P_2_2, a[2], b[2]);
	and A_2_3(P_2_3, a[2], b[3]);
	and A_2_4(P_2_4, a[2], b[4]);
	and A_2_5(P_2_5, a[2], b[5]);
	and A_2_6(P_2_6, a[2], b[6]);
	and A_2_7(P_2_7, a[2], b[7]);
	and A_2_8(P_2_8, a[2], b[8]);
	and A_2_9(P_2_9, a[2], b[9]);
	and A_2_10(P_2_10, a[2], b[10]);
	and A_2_11(P_2_11, a[2], b[11]);
	and A_2_12(P_2_12, a[2], b[12]);
	and A_2_13(P_2_13, a[2], b[13]);
	and A_2_14(P_2_14, a[2], b[14]);
	and A_2_15(P_2_15, a[2], b[15]);
	and A_3_0(P_3_0, a[3], b[0]);
	and A_3_1(P_3_1, a[3], b[1]);
	and A_3_2(P_3_2, a[3], b[2]);
	and A_3_3(P_3_3, a[3], b[3]);
	and A_3_4(P_3_4, a[3], b[4]);
	and A_3_5(P_3_5, a[3], b[5]);
	and A_3_6(P_3_6, a[3], b[6]);
	and A_3_7(P_3_7, a[3], b[7]);
	and A_3_8(P_3_8, a[3], b[8]);
	and A_3_9(P_3_9, a[3], b[9]);
	and A_3_10(P_3_10, a[3], b[10]);
	and A_3_11(P_3_11, a[3], b[11]);
	and A_3_12(P_3_12, a[3], b[12]);
	and A_3_13(P_3_13, a[3], b[13]);
	and A_3_14(P_3_14, a[3], b[14]);
	and A_3_15(P_3_15, a[3], b[15]);
	and A_4_0(P_4_0, a[4], b[0]);
	and A_4_1(P_4_1, a[4], b[1]);
	and A_4_2(P_4_2, a[4], b[2]);
	and A_4_3(P_4_3, a[4], b[3]);
	and A_4_4(P_4_4, a[4], b[4]);
	and A_4_5(P_4_5, a[4], b[5]);
	and A_4_6(P_4_6, a[4], b[6]);
	and A_4_7(P_4_7, a[4], b[7]);
	and A_4_8(P_4_8, a[4], b[8]);
	and A_4_9(P_4_9, a[4], b[9]);
	and A_4_10(P_4_10, a[4], b[10]);
	and A_4_11(P_4_11, a[4], b[11]);
	and A_4_12(P_4_12, a[4], b[12]);
	and A_4_13(P_4_13, a[4], b[13]);
	and A_4_14(P_4_14, a[4], b[14]);
	and A_4_15(P_4_15, a[4], b[15]);
	and A_5_0(P_5_0, a[5], b[0]);
	and A_5_1(P_5_1, a[5], b[1]);
	and A_5_2(P_5_2, a[5], b[2]);
	and A_5_3(P_5_3, a[5], b[3]);
	and A_5_4(P_5_4, a[5], b[4]);
	and A_5_5(P_5_5, a[5], b[5]);
	and A_5_6(P_5_6, a[5], b[6]);
	and A_5_7(P_5_7, a[5], b[7]);
	and A_5_8(P_5_8, a[5], b[8]);
	and A_5_9(P_5_9, a[5], b[9]);
	and A_5_10(P_5_10, a[5], b[10]);
	and A_5_11(P_5_11, a[5], b[11]);
	and A_5_12(P_5_12, a[5], b[12]);
	and A_5_13(P_5_13, a[5], b[13]);
	and A_5_14(P_5_14, a[5], b[14]);
	and A_5_15(P_5_15, a[5], b[15]);
	and A_6_0(P_6_0, a[6], b[0]);
	and A_6_1(P_6_1, a[6], b[1]);
	and A_6_2(P_6_2, a[6], b[2]);
	and A_6_3(P_6_3, a[6], b[3]);
	and A_6_4(P_6_4, a[6], b[4]);
	and A_6_5(P_6_5, a[6], b[5]);
	and A_6_6(P_6_6, a[6], b[6]);
	and A_6_7(P_6_7, a[6], b[7]);
	and A_6_8(P_6_8, a[6], b[8]);
	and A_6_9(P_6_9, a[6], b[9]);
	and A_6_10(P_6_10, a[6], b[10]);
	and A_6_11(P_6_11, a[6], b[11]);
	and A_6_12(P_6_12, a[6], b[12]);
	and A_6_13(P_6_13, a[6], b[13]);
	and A_6_14(P_6_14, a[6], b[14]);
	and A_6_15(P_6_15, a[6], b[15]);
	and A_7_0(P_7_0, a[7], b[0]);
	and A_7_1(P_7_1, a[7], b[1]);
	and A_7_2(P_7_2, a[7], b[2]);
	and A_7_3(P_7_3, a[7], b[3]);
	and A_7_4(P_7_4, a[7], b[4]);
	and A_7_5(P_7_5, a[7], b[5]);
	and A_7_6(P_7_6, a[7], b[6]);
	and A_7_7(P_7_7, a[7], b[7]);
	and A_7_8(P_7_8, a[7], b[8]);
	and A_7_9(P_7_9, a[7], b[9]);
	and A_7_10(P_7_10, a[7], b[10]);
	and A_7_11(P_7_11, a[7], b[11]);
	and A_7_12(P_7_12, a[7], b[12]);
	and A_7_13(P_7_13, a[7], b[13]);
	and A_7_14(P_7_14, a[7], b[14]);
	and A_7_15(P_7_15, a[7], b[15]);
	and A_8_0(P_8_0, a[8], b[0]);
	and A_8_1(P_8_1, a[8], b[1]);
	and A_8_2(P_8_2, a[8], b[2]);
	and A_8_3(P_8_3, a[8], b[3]);
	and A_8_4(P_8_4, a[8], b[4]);
	and A_8_5(P_8_5, a[8], b[5]);
	and A_8_6(P_8_6, a[8], b[6]);
	and A_8_7(P_8_7, a[8], b[7]);
	and A_8_8(P_8_8, a[8], b[8]);
	and A_8_9(P_8_9, a[8], b[9]);
	and A_8_10(P_8_10, a[8], b[10]);
	and A_8_11(P_8_11, a[8], b[11]);
	and A_8_12(P_8_12, a[8], b[12]);
	and A_8_13(P_8_13, a[8], b[13]);
	and A_8_14(P_8_14, a[8], b[14]);
	and A_8_15(P_8_15, a[8], b[15]);
	and A_9_0(P_9_0, a[9], b[0]);
	and A_9_1(P_9_1, a[9], b[1]);
	and A_9_2(P_9_2, a[9], b[2]);
	and A_9_3(P_9_3, a[9], b[3]);
	and A_9_4(P_9_4, a[9], b[4]);
	and A_9_5(P_9_5, a[9], b[5]);
	and A_9_6(P_9_6, a[9], b[6]);
	and A_9_7(P_9_7, a[9], b[7]);
	and A_9_8(P_9_8, a[9], b[8]);
	and A_9_9(P_9_9, a[9], b[9]);
	and A_9_10(P_9_10, a[9], b[10]);
	and A_9_11(P_9_11, a[9], b[11]);
	and A_9_12(P_9_12, a[9], b[12]);
	and A_9_13(P_9_13, a[9], b[13]);
	and A_9_14(P_9_14, a[9], b[14]);
	and A_9_15(P_9_15, a[9], b[15]);
	and A_10_0(P_10_0, a[10], b[0]);
	and A_10_1(P_10_1, a[10], b[1]);
	and A_10_2(P_10_2, a[10], b[2]);
	and A_10_3(P_10_3, a[10], b[3]);
	and A_10_4(P_10_4, a[10], b[4]);
	and A_10_5(P_10_5, a[10], b[5]);
	and A_10_6(P_10_6, a[10], b[6]);
	and A_10_7(P_10_7, a[10], b[7]);
	and A_10_8(P_10_8, a[10], b[8]);
	and A_10_9(P_10_9, a[10], b[9]);
	and A_10_10(P_10_10, a[10], b[10]);
	and A_10_11(P_10_11, a[10], b[11]);
	and A_10_12(P_10_12, a[10], b[12]);
	and A_10_13(P_10_13, a[10], b[13]);
	and A_10_14(P_10_14, a[10], b[14]);
	and A_10_15(P_10_15, a[10], b[15]);
	and A_11_0(P_11_0, a[11], b[0]);
	and A_11_1(P_11_1, a[11], b[1]);
	and A_11_2(P_11_2, a[11], b[2]);
	and A_11_3(P_11_3, a[11], b[3]);
	and A_11_4(P_11_4, a[11], b[4]);
	and A_11_5(P_11_5, a[11], b[5]);
	and A_11_6(P_11_6, a[11], b[6]);
	and A_11_7(P_11_7, a[11], b[7]);
	and A_11_8(P_11_8, a[11], b[8]);
	and A_11_9(P_11_9, a[11], b[9]);
	and A_11_10(P_11_10, a[11], b[10]);
	and A_11_11(P_11_11, a[11], b[11]);
	and A_11_12(P_11_12, a[11], b[12]);
	and A_11_13(P_11_13, a[11], b[13]);
	and A_11_14(P_11_14, a[11], b[14]);
	and A_11_15(P_11_15, a[11], b[15]);
	and A_12_0(P_12_0, a[12], b[0]);
	and A_12_1(P_12_1, a[12], b[1]);
	and A_12_2(P_12_2, a[12], b[2]);
	and A_12_3(P_12_3, a[12], b[3]);
	and A_12_4(P_12_4, a[12], b[4]);
	and A_12_5(P_12_5, a[12], b[5]);
	and A_12_6(P_12_6, a[12], b[6]);
	and A_12_7(P_12_7, a[12], b[7]);
	and A_12_8(P_12_8, a[12], b[8]);
	and A_12_9(P_12_9, a[12], b[9]);
	and A_12_10(P_12_10, a[12], b[10]);
	and A_12_11(P_12_11, a[12], b[11]);
	and A_12_12(P_12_12, a[12], b[12]);
	and A_12_13(P_12_13, a[12], b[13]);
	and A_12_14(P_12_14, a[12], b[14]);
	and A_12_15(P_12_15, a[12], b[15]);
	and A_13_0(P_13_0, a[13], b[0]);
	and A_13_1(P_13_1, a[13], b[1]);
	and A_13_2(P_13_2, a[13], b[2]);
	and A_13_3(P_13_3, a[13], b[3]);
	and A_13_4(P_13_4, a[13], b[4]);
	and A_13_5(P_13_5, a[13], b[5]);
	and A_13_6(P_13_6, a[13], b[6]);
	and A_13_7(P_13_7, a[13], b[7]);
	and A_13_8(P_13_8, a[13], b[8]);
	and A_13_9(P_13_9, a[13], b[9]);
	and A_13_10(P_13_10, a[13], b[10]);
	and A_13_11(P_13_11, a[13], b[11]);
	and A_13_12(P_13_12, a[13], b[12]);
	and A_13_13(P_13_13, a[13], b[13]);
	and A_13_14(P_13_14, a[13], b[14]);
	and A_13_15(P_13_15, a[13], b[15]);
	and A_14_0(P_14_0, a[14], b[0]);
	and A_14_1(P_14_1, a[14], b[1]);
	and A_14_2(P_14_2, a[14], b[2]);
	and A_14_3(P_14_3, a[14], b[3]);
	and A_14_4(P_14_4, a[14], b[4]);
	and A_14_5(P_14_5, a[14], b[5]);
	and A_14_6(P_14_6, a[14], b[6]);
	and A_14_7(P_14_7, a[14], b[7]);
	and A_14_8(P_14_8, a[14], b[8]);
	and A_14_9(P_14_9, a[14], b[9]);
	and A_14_10(P_14_10, a[14], b[10]);
	and A_14_11(P_14_11, a[14], b[11]);
	and A_14_12(P_14_12, a[14], b[12]);
	and A_14_13(P_14_13, a[14], b[13]);
	and A_14_14(P_14_14, a[14], b[14]);
	and A_14_15(P_14_15, a[14], b[15]);
	and A_15_0(P_15_0, a[15], b[0]);
	and A_15_1(P_15_1, a[15], b[1]);
	and A_15_2(P_15_2, a[15], b[2]);
	and A_15_3(P_15_3, a[15], b[3]);
	and A_15_4(P_15_4, a[15], b[4]);
	and A_15_5(P_15_5, a[15], b[5]);
	and A_15_6(P_15_6, a[15], b[6]);
	and A_15_7(P_15_7, a[15], b[7]);
	and A_15_8(P_15_8, a[15], b[8]);
	and A_15_9(P_15_9, a[15], b[9]);
	and A_15_10(P_15_10, a[15], b[10]);
	and A_15_11(P_15_11, a[15], b[11]);
	and A_15_12(P_15_12, a[15], b[12]);
	and A_15_13(P_15_13, a[15], b[13]);
	and A_15_14(P_15_14, a[15], b[14]);
	and A_15_15(P_15_15, a[15], b[15]);
	//-------------------------------------------layer 1---------------------------------------//  
	wire SH_1;
	wire SH_2;
	wire SH_3;
	wire SH_4;
 	
	wire CH_1;
	wire CH_2;
	wire CH_3;
	wire CH_4;

	wire SF_1;
	wire SF_2;
	wire SF_3;
	wire SF_4;
	wire SF_5;
	wire SF_6;
	wire SF_7;
	wire SF_8;
 	
	wire CF_1;
	wire CF_2;
	wire CF_3;
	wire CF_4;
	wire CF_5;
	wire CF_6;
	wire CF_7;
	wire CF_8;

	wire SC_1;
	wire SC_2;
	wire SC_3;
	wire SC_4;
	wire SC_5;
	wire SC_6;
	wire SC_7;
	wire SC_8;
	wire SC_9;
	wire SC_10;
	wire SC_11;
	wire SC_12;
	wire SC_13;
	wire SC_14;
	wire SC_15;
	wire SC_16;
	wire SC_17;
	wire SC_18;
	wire SC_19;
	wire SC_20;
	wire SC_21;
	wire SC_22;
	wire SC_23;
	wire SC_24;
	wire SC_25;
	wire SC_26;
	wire SC_27;
	wire SC_28;
	wire SC_29;
	wire SC_30;
	wire SC_31;
	wire SC_32;
	wire SC_33;
	wire SC_34;
	wire SC_35;
	wire SC_36;
	wire SC_37;
	wire SC_38;
	wire SC_39;
	wire SC_40;
	wire SC_41;
	wire SC_42;
	wire SC_43;
	wire SC_44;
	wire SC_45;
	wire SC_46;
	wire SC_47;
	wire SC_48;
	wire SC_49;
	wire SC_50;
	wire SC_51;
	wire SC_52;
	wire SC_53;
	wire SC_54;
	wire SC_55;
	wire SC_56;

	wire CC_1;
	wire CC_2;
	wire CC_3;
	wire CC_4;
	wire CC_5;
	wire CC_6;
	wire CC_7;
	wire CC_8;
	wire CC_9;
	wire CC_10;
	wire CC_11;
	wire CC_12;
	wire CC_13;
	wire CC_14;
	wire CC_15;
	wire CC_16;
	wire CC_17;
	wire CC_18;
	wire CC_19;
	wire CC_20;
	wire CC_21;
	wire CC_22;
	wire CC_23;
	wire CC_24;
	wire CC_25;
	wire CC_26;
	wire CC_27;
	wire CC_28;
	wire CC_29;
	wire CC_30;
	wire CC_31;
	wire CC_32;
	wire CC_33;
	wire CC_34;
	wire CC_35;
	wire CC_36;
	wire CC_37;
	wire CC_38;
	wire CC_39;
	wire CC_40;
	wire CC_41;
	wire CC_42;
	wire CC_43;
	wire CC_44;
	wire CC_45;
	wire CC_46;
	wire CC_47;
	wire CC_48;
	wire CC_49;
	wire CC_50;
	wire CC_51;
	wire CC_52;
	wire CC_53;
	wire CC_54;
	wire CC_55;
	wire CC_56;
 	
	wire CO_1;
	wire CO_2;
	wire CO_3;
	wire CO_4;
	wire CO_5;
	wire CO_6;
	wire CO_7;
	wire CO_8;
	wire CO_9;
	wire CO_10;
	wire CO_11;
	wire CO_12;
	wire CO_13;
	wire CO_14;
	wire CO_15;
	wire CO_16;
	wire CO_17;
	wire CO_18;
	wire CO_19;
	wire CO_20;
	wire CO_21;
	wire CO_22;
	wire CO_23;
	wire CO_24;
	wire CO_25;
	wire CO_26;
	wire CO_27;
	wire CO_28;
	wire CO_29;
	wire CO_30;
	wire CO_31;
	wire CO_32;
	wire CO_33;
	wire CO_34;
	wire CO_35;
	wire CO_36;
	wire CO_37;
	wire CO_38;
	wire CO_39;
	wire CO_40;
	wire CO_41;
	wire CO_42;
	wire CO_43;
	wire CO_44;
	wire CO_45;
	wire CO_46;
	wire CO_47;
	wire CO_48;
	wire CO_49;
	wire CO_50;
	wire CO_51;
	wire CO_52;
	wire CO_53;
	wire CO_54;
	wire CO_55;
	wire CO_56;

	//half adder
	ha HA_1(SH_1, CH_1, P_0_1, P_1_0);
	ha HA_2(SH_2, CH_2, P_1_4, P_0_5);
	ha HA_3(SH_3, CH_3, P_1_8, P_0_9);
	ha HA_4(SH_4, CH_4, P_1_12, P_0_13);
 	
	//full adder
	fa FA_1(SF_1, CF_1, P_2_0, P_1_1, P_0_2);
	fa FA_2(SF_2, CF_2, P_15_2, P_14_3, CO_14);
	fa FA_3(SF_3, CF_3, P_2_4, P_1_5, P_0_6);
	fa FA_4(SF_4, CF_4, P_15_6, P_14_7, CO_28);
	fa FA_5(SF_5, CF_5, P_2_8, P_1_9, P_0_10);
	fa FA_6(SF_6, CF_6, P_15_10, P_14_11, CO_42);
	fa FA_7(SF_7, CF_7, P_2_12, P_1_13, P_0_4);
	fa FA_8(SF_8, CF_8, P_15_14, P_14_15, CO_56);
 	
	//compressor;
	cp_acc CP_1(SC_1,CO_1,CC_1,P_3_0,P_2_1,P_1_2,P_0_3,ground_z);
	cp_acc CP_2(SC_2,CO_2,CC_2,P_4_0,P_3_1,P_2_2,P_1_3,CO_1);
	cp_acc CP_3(SC_3,CO_3,CC_3,P_5_0,P_4_1,P_3_2,P_2_3,CO_2);
	cp_acc CP_4(SC_4,CO_4,CC_4,P_6_0,P_5_1,P_4_2,P_3_3,CO_3);
	cp_acc CP_5(SC_5,CO_5,CC_5,P_7_0,P_6_1,P_5_2,P_4_2,CO_4);
	cp_acc CP_6(SC_6,CO_6,CC_6,P_8_0,P_7_1,P_6_2,P_5_3,CO_5);
	cp_acc CP_7(SC_7,CO_7,CC_7,P_9_0,P_8_1,P_7_2,P_6_3,CO_6);
	cp_acc CP_8(SC_8,CO_8,CC_8,P_10_0,P_9_1,P_8_2,P_7_3,CO_7);
	cp_acc CP_9(SC_9,CO_9,CC_9,P_11_0,P_10_1,P_9_2,P_8_3,CO_8);
	cp_acc CP_10(SC_10,CO_10,CC_10,P_12_0,P_11_1,P_10_2,P_9_3,CO_9);
	cp_acc CP_11(SC_11,CO_11,CC_11,P_13_0,P_12_1,P_11_2,P_10_3,CO_10);
	cp_acc CP_12(SC_12,CO_12,CC_12,P_14_0,P_13_1,P_12_2,P_11_3,CO_11);
	cp_acc CP_13(SC_13,CO_13,CC_13,P_15_0,P_14_1,P_13_2,P_12_3,CO_12);
	cp_acc CP_14(SC_14,CO_14,CC_14,P_15_1,P_14_2,P_13_3,ground_z,CO_13);
	cp_acc CP_15(SC_15,CO_15,CC_15,P_3_4,P_2_5,P_1_6,P_0_7,ground_z);
	cp_acc CP_16(SC_16,CO_16,CC_16,P_4_4,P_3_5,P_2_6,P_1_7,CO_15);
	cp_acc CP_17(SC_17,CO_17,CC_17,P_5_4,P_4_5,P_3_6,P_2_7,CO_16);
	cp_acc CP_18(SC_18,CO_18,CC_18,P_6_4,P_5_5,P_4_6,P_3_7,CO_17);
	cp_acc CP_19(SC_19,CO_19,CC_19,P_7_4,P_6_5,P_5_6,P_4_7,CO_18);
	cp_acc CP_20(SC_20,CO_20,CC_20,P_8_4,P_7_5,P_6_6,P_5_7,CO_19);
	cp_acc CP_21(SC_21,CO_21,CC_21,P_9_4,P_8_5,P_7_6,P_6_7,CO_20);
	cp_acc CP_22(SC_22,CO_22,CC_22,P_10_4,P_9_5,P_8_6,P_7_7,CO_21);
	cp_acc CP_23(SC_23,CO_23,CC_23,P_11_4,P_10_5,P_9_6,P_8_7,CO_22);
	cp_acc CP_24(SC_24,CO_24,CC_24,P_12_4,P_11_5,P_10_6,P_9_7,CO_23);
	cp_acc CP_25(SC_25,CO_25,CC_25,P_13_4,P_12_5,P_11_6,P_10_7,CO_24);
	cp_acc CP_26(SC_26,CO_26,CC_26,P_14_4,P_13_5,P_12_6,P_11_7,CO_25);
	cp_acc CP_27(SC_27,CO_27,CC_27,P_15_4,P_14_5,P_13_6,P_12_7,CO_26);
	cp_acc CP_28(SC_28,CO_28,CC_28,P_15_4,P_14_6,P_13_7,ground_z,CO_27);
	cp_acc CP_29(SC_29,CO_29,CC_29,P_3_8,P_2_9,P_1_10,P_0_11,ground_z);
	cp_acc CP_30(SC_30,CO_30,CC_30,P_4_8,P_3_9,P_2_10,P_1_11,CO_29);
	cp_acc CP_31(SC_31,CO_31,CC_31,P_5_8,P_4_9,P_3_10,P_2_11,CO_30);
	cp_acc CP_32(SC_32,CO_32,CC_32,P_6_8,P_5_9,P_4_10,P_3_11,CO_31);
	cp_acc CP_33(SC_33,CO_33,CC_33,P_7_8,P_6_9,P_5_10,P_4_11,CO_32);
	cp_acc CP_34(SC_34,CO_34,CC_34,P_8_8,P_7_9,P_6_10,P_5_11,CO_33);
	cp_acc CP_35(SC_35,CO_35,CC_35,P_9_8,P_8_9,P_7_10,P_6_11,CO_34);
	cp_acc CP_36(SC_36,CO_36,CC_36,P_10_8,P_9_9,P_8_10,P_7_11,CO_35);
	cp_acc CP_37(SC_37,CO_37,CC_37,P_11_8,P_10_9,P_9_10,P_8_11,CO_36);
	cp_acc CP_38(SC_38,CO_38,CC_38,P_12_8,P_11_9,P_10_10,P_9_11,CO_37);
	cp_acc CP_39(SC_39,CO_39,CC_39,P_13_8,P_12_9,P_11_10,P_10_11,CO_38);
	cp_acc CP_40(SC_40,CO_40,CC_40,P_14_8,P_13_9,P_12_10,P_11_11,CO_39);
	cp_acc CP_41(SC_41,CO_41,CC_41,P_15_8,P_14_9,P_13_10,P_12_11,CO_40);
	cp_acc CP_42(SC_42,CO_42,CC_42,P_15_9,P_14_10,P_13_11,ground_z,CO_41);
	cp_acc CP_43(SC_43,CO_43,CC_43,P_3_12,P_2_13,P_1_14,P_0_15,ground_z);
	cp_acc CP_44(SC_44,CO_44,CC_44,P_4_12,P_3_13,P_2_14,P_1_15,CO_43);
	cp_acc CP_45(SC_45,CO_45,CC_45,P_5_12,P_4_13,P_3_14,P_2_15,CO_44);
	cp_acc CP_46(SC_46,CO_46,CC_46,P_6_12,P_5_13,P_4_14,P_3_15,CO_45);
	cp_acc CP_47(SC_47,CO_47,CC_47,P_7_12,P_6_13,P_5_14,P_4_15,CO_46);
	cp_acc CP_48(SC_48,CO_48,CC_48,P_8_12,P_7_13,P_6_14,P_5_15,CO_47);
	cp_acc CP_49(SC_49,CO_49,CC_49,P_9_12,P_8_13,P_7_14,P_6_15,CO_48);
	cp_acc CP_50(SC_50,CO_50,CC_50,P_10_12,P_9_13,P_8_14,P_7_15,CO_49);
	cp_acc CP_51(SC_51,CO_51,CC_51,P_11_12,P_10_13,P_9_14,P_8_15,CO_50);
	cp_acc CP_52(SC_52,CO_52,CC_52,P_12_12,P_11_13,P_10_14,P_9_15,CO_51);
	cp_acc CP_53(SC_53,CO_53,CC_53,P_13_12,P_12_13,P_11_14,P_10_15,CO_52);
	cp_acc CP_54(SC_54,CO_54,CC_54,P_14_12,P_13_13,P_12_14,P_11_15,CO_53);
	cp_acc CP_55(SC_55,CO_55,CC_55,P_15_12,P_14_13,P_13_14,P_12_15,CO_54);
	cp_acc CP_56(SC_56,CO_56,CC_56,P_15_13,P_14_14,P_13_15,ground_z,CO_55);

	//-------------------------------------------layer 2---------------------------------------//  
	wire SH_5;
	wire SH_6;
	wire SH_7;
	wire SH_8;
	wire SH_9;
	wire SH_10;
	wire SH_11;
	wire SH_12;
	wire SH_13;
	wire SH_14;
 	
	wire CH_5;
	wire CH_6;
	wire CH_7;
	wire CH_8;
	wire CH_9;
	wire CH_10;
	wire CH_11;
	wire CH_12;
	wire CH_13;
	wire CH_14;

	wire SF_9;
	wire SF_10;
	wire SF_11;
	wire SF_12;
	wire SF_13;
	wire SF_14;

	wire CF_9;
	wire CF_10;
	wire CF_11;
	wire CF_12;
	wire CF_13;
	wire CF_14;
 	
	wire SC_57;
	wire SC_58;
	wire SC_59;
	wire SC_60;
	wire SC_61;
	wire SC_62;
	wire SC_63;
	wire SC_64;
	wire SC_65;
	wire SC_66;
	wire SC_67;
	wire SC_68;
	wire SC_69;
	wire SC_70;
	wire SC_71;
	//wire SC_72;
	wire SC_73;
	wire SC_74;
	wire SC_75;
	wire SC_76;
	wire SC_77;
	wire SC_78;
	wire SC_79;
	wire SC_80;
	wire SC_81;
	wire SC_82;
	wire SC_83;

	wire CC_57;
	wire CC_58;
	wire CC_59;
	wire CC_60;
	wire CC_61;
	wire CC_62;
	wire CC_63;
	wire CC_64;
	wire CC_65;
	wire CC_66;
	wire CC_67;
	wire CC_68;
	wire CC_69;
	wire CC_70;
	wire CC_71;
	//wire CC_72;
	wire CC_73;
	wire CC_74;
	wire CC_75;
	wire CC_76;
	wire CC_77;
	wire CC_78;
	wire CC_79;
	wire CC_80;
	wire CC_81;
	wire CC_82;
	wire CC_83;

	wire CO_57;
	wire CO_58;
	wire CO_59;
	wire CO_60;
	wire CO_61;
	wire CO_62;
	wire CO_63;
	wire CO_64;
	wire CO_65;
	wire CO_66;
	wire CO_67;
	wire CO_68;
	wire CO_69;
	wire CO_70;
	wire CO_71;
	//wire CO_72;
	wire CO_73;
	wire CO_74;
	wire CO_75;
	wire CO_76;
	wire CO_77;
	wire CO_78;
	wire CO_79;
	wire CO_80;
	wire CO_81;
	wire CO_82;
	wire CO_83;

	
	//half adder
 	
	ha HA_5(SH_5, CH_5, SF_1, CH_1);
	ha HA_6(SH_6, CH_6, SC_1, CF_1);
	ha HA_7(SH_7, CH_7, SC_28, CC_27);
	ha HA_8(SH_8, CH_8, SF_4, CC_28);
	ha HA_9(SH_9, CH_9, CF_4, P_15_7);
	ha HA_10(SH_10, CH_10, SF_5, CH_3);
	ha HA_11(SH_11, CH_11, SC_29, CF_5);
	ha HA_12(SH_12, CH_12, SC_56, CC_54);
	ha HA_13(SH_13, CH_13, SC_56, CC_56);
	ha HA_14(SH_14, CH_14, CF_8, P_15_15);
 	
	//full adder
	fa FA_9(SF_9, CF_9, SC_2, CC_1, P_0_4);
	fa FA_10(SF_10, CF_10, SC_3, CC_2, SH_2);
	fa FA_11(SF_11, CF_11, SC_27, CC_26, CO_69);
	fa FA_12(SF_12, CF_12, SC_30, CC_29, P_0_12);
	fa FA_13(SF_13, CF_13, SC_31, CC_30, SH_4);
	fa FA_14(SF_14, CF_14, SC_55, CC_54, CO_83);
 	
 	
	//compressor
	cp_acc CP_57(SC_57,CO_57,CC_57,SC_4,CC_3,SF_3,CH_2,ground_z);
	cp_acc CP_58(SC_58,CO_58,CC_58,SC_5,CC_4,SC_15,CF_3,CO_57);
	cp_acc CP_59(SC_59,CO_59,CC_59,SC_6,CC_5,SC_16,CC_15,CO_58);
	cp_acc CP_60(SC_60,CO_60,CC_60,SC_7,CC_6,SC_17,CC_16,CO_59);
	cp_acc CP_61(SC_61,CO_61,CC_61,SC_8,CC_7,SC_18,CC_17,CO_60);
	cp_acc CP_62(SC_62,CO_62,CC_62,SC_9,CC_8,SC_19,CC_18,CO_61);
	cp_acc CP_63(SC_63,CO_63,CC_63,SC_10,CC_9,SC_20,CC_19,CO_62);
	cp_acc CP_64(SC_64,CO_64,CC_64,SC_11,CC_10,SC_21,CC_20,CO_63);
	cp_acc CP_65(SC_65,CO_65,CC_65,SC_12,CC_11,SC_22,CC_21,CO_64);
	cp_acc CP_66(SC_66,CO_66,CC_66,SC_13,CC_12,SC_23,CC_22,CO_65);
	cp_acc CP_67(SC_67,CO_67,CC_67,SC_14,CC_13,SC_24,CC_23,CO_66);
	cp_acc CP_68(SC_68,CO_68,CC_68,SF_2,CC_14,SC_25,CC_24,CO_67);
	cp_acc CP_69(SC_69,CO_69,CC_69,CF_2,P_15_3,SC_26,CC_25,CO_68);
	cp_acc CP_70(SC_70,CO_70,CC_70,SC_32,CC_31,SF_7,CH_4,ground_z);
	cp_acc CP_71(SC_71,CO_71,CC_71,SC_33,CC_32,SC_43,CF_7,CO_70);
	//cp_a CP_72cc(SC_72,CO_72,CC_72,SC_34,CC_44,SC_15,CF_3,CO_57);
	cp_acc CP_73(SC_73,CO_73,CC_73,SC_34,CC_33,SC_44,CC_43,CO_71);
	cp_acc CP_74(SC_74,CO_74,CC_74,SC_35,CC_34,SC_45,CC_44,CO_73);
	cp_acc CP_75(SC_75,CO_75,CC_75,SC_36,CC_35,SC_46,CC_45,CO_74);
	cp_acc CP_76(SC_76,CO_76,CC_76,SC_37,CC_36,SC_47,CC_46,CO_75);
	cp_acc CP_77(SC_77,CO_77,CC_77,SC_38,CC_37,SC_48,CC_47,CO_76);
	cp_acc CP_78(SC_78,CO_78,CC_78,SC_39,CC_38,SC_49,CC_48,CO_77);
	cp_acc CP_79(SC_79,CO_79,CC_79,SC_40,CC_39,SC_50,CC_49,CO_78);
	cp_acc CP_80(SC_80,CO_80,CC_80,SC_41,CC_40,SC_51,CC_50,CO_79);
	cp_acc CP_81(SC_81,CO_81,CC_81,SC_42,CC_41,SC_52,CC_51,CO_80);
	cp_acc CP_82(SC_82,CO_82,CC_82,SF_6,CC_42,SC_53,CC_52,CO_81);
	cp_acc CP_83(SC_83,CO_83,CC_83,CF_6,P_15_11,SC_54,CC_53,CO_82);

 	
	//-------------------------------------------layer 3---------------------------------------//  ;
	wire SH_15;
	wire SH_16;
	wire SH_17;
	wire SH_18;
	wire SH_19;
	wire SH_20;
	wire SH_21;
	wire SH_22;
	wire SH_23;
	wire SH_24;
	wire SH_25;
 	

	wire CH_15;
	wire CH_16;
	wire CH_17;
	wire CH_18;
	wire CH_19;
	wire CH_20;
	wire CH_21;
	wire CH_22;
	wire CH_23;
	wire CH_24;
	wire CH_25;

	wire SF_15;
	wire SF_16;
	wire SF_17;
	wire SF_18;
 	
	wire CF_15;
	wire CF_16;
	wire CF_17;
	wire CF_18;

	wire SC_84;
	wire SC_85;
	wire SC_86;
	wire SC_87;
	wire SC_88;
	wire SC_89;
	wire SC_90;
	wire SC_91;
	wire SC_92;
	wire SC_93;
	wire SC_94;
	wire SC_95;
	wire SC_96;

	wire CC_84;
	wire CC_85;
	wire CC_86;
	wire CC_87;
	wire CC_88;
	wire CC_89;
	wire CC_90;
	wire CC_91;
	wire CC_92;
	wire CC_93;
	wire CC_94;
	wire CC_95;
	wire CC_96;

	wire CO_84;
	wire CO_85;
	wire CO_86;
	wire CO_87;
	wire CO_88;
	wire CO_89;
	wire CO_90;
	wire CO_91;
	wire CO_92;
	wire CO_93;
	wire CO_94;
	wire CO_95;
	wire CO_96;

	
	//half adder
 	
	ha HA_15(SH_15, CH_15, SH_6, CH_5);
	ha HA_16(SH_16, CH_16, SF_9, CH_6);
	ha HA_17(SH_17, CH_17, SF_10, CF_9);
	ha HA_18(SH_18, CH_18, SC_57, CF_10);
	ha HA_19(SH_19, CH_19, SC_58, CC_57);
	ha HA_20(SH_20, CH_20, SC_82, CC_81);
	ha HA_21(SH_21, CH_21, SC_83, CC_82);
	ha HA_22(SH_22, CH_22, SF_14, CC_83);
	ha HA_23(SH_23, CH_23, SH_12, CF_14);
	ha HA_24(SH_24, CH_24, SH_13, CH_12);
	ha HA_25(SH_25, CH_25, SH_14, CH_13);
 	
	//full adder
	fa FA_15(SF_15, CF_15, SC_59, CC_58, P_0_8);
	fa FA_16(SF_16, CF_16, SC_60, CC_59, SH_3);
	fa FA_17(SF_17, CF_17, SC_61, CC_60, SH_10);
	fa FA_18(SF_18, CF_18, SC_81, CC_80, CO_96);
 	
	cp_acc CP_84(SC_84,CO_84,CC_84,SC_62,CC_61,SH_11,CH_10,ground_z);
	cp_acc CP_85(SC_85,CO_85,CC_85,SC_63,CC_62,SH_12,CH_11,CO_84);
	cp_acc CP_86(SC_86,CO_86,CC_86,SC_64,CC_63,SH_13,CH_12,CO_85);
	cp_acc CP_87(SC_87,CO_87,CC_87,SC_65,CC_64,SC_70,CH_13,CO_86);
	cp_acc CP_88(SC_88,CO_88,CC_88,SC_66,CC_65,SC_71,CC_70,CO_87);
	cp_acc CP_89(SC_89,CO_89,CC_89,SC_67,CC_66,SC_73,CC_71,CO_88);
	cp_acc CP_90(SC_90,CO_90,CC_90,SC_68,CC_67,SC_74,CC_73,CO_89);
	cp_acc CP_91(SC_91,CO_91,CC_91,SC_69,CC_68,SC_75,CC_74,CO_90);
	cp_acc CP_92(SC_92,CO_92,CC_92,SF_11,CC_69,SC_76,CC_75,CO_91);
	cp_acc CP_93(SC_93,CO_93,CC_93,SH_7,CF_11,SC_77,CC_76,CO_92);
	cp_acc CP_94(SC_94,CO_94,CC_94,SH_8,CH_7,SC_78,CC_77,CO_93);
	cp_acc CP_95(SC_95,CO_95,CC_95,SH_9,CH_8,SC_79,CC_78,CO_94);
	cp_acc CP_96(SC_96,CO_96,CC_96,CH_9,SC_80,CC_79,ground_z,CO_95);
 	
 	
	//results
	wire CF_26;
	wire CF_27;
	wire CF_28;
	wire CF_29;
	wire CF_30;
	wire CF_31;
	wire CF_32;
	wire CF_33;
	wire CF_34;
	wire CF_35;
	wire CF_36;
	wire CF_37;
	wire CF_38;
	wire CF_39;
	wire CF_40;
	wire CF_41;
	wire CF_42;
	wire CF_43;
	wire CF_44;
	wire CF_45;
	wire CF_46;
	wire CF_47;
	wire CF_48;
	wire CF_49;
	wire CF_50;
	wire CF_51;
	wire CF_52;
  
	wire SF_26;
	wire SF_27;
	wire SF_28;
	wire SF_29;
	wire SF_30;
	wire SF_31;
	wire SF_32;
	wire SF_33;
	wire SF_34;
	wire SF_35;
	wire SF_36;
	wire SF_37;
	wire SF_38;
	wire SF_39;
	wire SF_40;
	wire SF_41;
	wire SF_42;
	wire SF_43;
	wire SF_44;
	wire SF_45;
	wire SF_46;
	wire SF_47;
	wire SF_48;
	wire SF_49;
	wire SF_50;
	wire SF_51;
	wire SF_52;

	fa FA_19(SF_26, CF_26, SH_16, CH_15,ground_z);
	fa FA_20(SF_27, CF_27, SH_17, CH_16,CF_26);
	fa FA_21(SF_28, CF_28, SH_18, CH_17,CF_27);
	fa FA_22(SF_29, CF_29, SH_19, CH_18,CF_28);
	fa FA_23(SF_30, CF_30, SF_15, CH_19,CF_29);
	fa FA_24(SF_31, CF_31, SF_16, CF_15,CF_30);
	fa FA_25(SF_32, CF_32, SF_17, CF_16,CF_31);
	fa FA_26(SF_33, CF_33, SC_84, CF_17,CF_32);
	fa FA_27(SF_34, CF_34, SC_85, CC_84,CF_33);
	fa FA_28(SF_35, CF_35, SC_86, CC_85,CF_34);
	fa FA_29(SF_36, CF_36, SC_87, CC_86,CF_35);
	fa FA_30(SF_37, CF_37, SC_88, CC_87,CF_36);
	fa FA_31(SF_38, CF_38, SC_89, CC_88,CF_37);
	fa FA_32(SF_39, CF_39, SC_90, CC_89,CF_38);
	fa FA_33(SF_40, CF_40, SC_91, CC_90,CF_39);
	fa FA_34(SF_41, CF_41, SC_92, CC_91,CF_40);
	fa FA_35(SF_42, CF_42, SC_93, CC_92,CF_41);
	fa FA_36(SF_43, CF_43, SC_94, CC_93,CF_42);
	fa FA_37(SF_44, CF_44, SC_95, CC_94,CF_43);
	fa FA_38(SF_45, CF_45, SC_96, CC_95,CF_44);
	fa FA_39(SF_46, CF_46, SF_18, CC_96,CF_45);
	fa FA_40(SF_47, CF_47, SH_20, CF_18,CF_46);
	fa FA_41(SF_48, CF_48, SH_21, CH_20,CF_47);
	fa FA_42(SF_49, CF_49, SH_22, CH_21,CF_48);
	fa FA_43(SF_50, CF_50, SH_23, CH_22,CF_49);
	fa FA_44(SF_51, CF_51, SH_24, CH_23,CF_50);
	fa FA_45(SF_52, CF_52, SH_25, CH_24,CF_51);
	fa FA_46(SF_53, CF_53, CH_25, CH_14,CF_52);
	assign sum = {SF_53,SF_52,SF_51,SF_50,SF_49,SF_48,SF_47,SF_46,SF_45,SF_44,SF_43,SF_42,SF_41,SF_40,SF_39,SF_38,SF_37,SF_36,SF_35,SF_34,SF_33,SF_32,SF_31,SF_30,SF_29,SF_28,SF_27,SF_26,SH_15,SH_5,SH_1,P_0_0};







	
endmodule


